package state_machine_pack is 
	
	type st is (st_0, st_1, st_2, st_3, st_4, st_5)
	
end state_machine_pack;